// module scoring_module (
// 	input clk,
// 	input reset,
// 	input ack,
// 	input bright,
//     input [9:0] pacX,
//     input [9:0] pacY,
// 	input [9:0] hCount, vCount,
// 	input [479:0] maze [639:0],
// 	input [479:0] intersection [639:0],
// 	input winIn,
// 	input loseIn,
// 	input [3:0] ghostFills,
// 	input pacmanFill,
// 	output reg [15:0] score,
// 	output reg [11:0] rgb,
// 	output winOut,
// 	output loseOut
//     );

// 	reg [4:0] state;
	
// 	localparam
// 	INI = 5'b00001;
// 	STANDBY = 5'b00010;
// 	WIN = 5'b00100;
// 	LOSE = 5'b01000;
	


// 	always@ (*) begin

// 	end













// endmodule